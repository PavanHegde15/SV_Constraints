module test();






endmodule
